module alu(
    input logic [2:0] control,
    input logic [31:0] input1,
    input logic [31:0] input2,
    output logic zero,
    output logic [31:0] result
);

    assign zero = result == 0;

    always_comb
        case(control)
            'b000: result = input1 + input2;
            'b001: result = input1 - input2;
            'b111: result = input1 & input2;
            default: $display("ALU: Control=0b%0b; Not handled", control);
        endcase

endmodule
